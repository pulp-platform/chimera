// Copyright 2024 ETH Zurich and University of Bologna.
// Solderpad Hardware License, Version 0.51, see LICENSE for details.
// SPDX-License-Identifier: SHL-0.51
//
// Moritz Scherer <scheremo@iis.ee.ethz.ch>

module chimera_cluster
  import chimera_pkg::*;
  import cheshire_pkg::*;
#(
  parameter cheshire_cfg_t Cfg = '0,

  parameter int unsigned NrCores           = 9,
  parameter type         narrow_in_req_t   = logic,
  parameter type         narrow_in_resp_t  = logic,
  parameter type         narrow_out_req_t  = logic,
  parameter type         narrow_out_resp_t = logic,
  parameter type         wide_out_req_t    = logic,
  parameter type         wide_out_resp_t   = logic,

  // !! DO NOT OVERWRITE THESE PARAMETERS
  // These parameters are used to provide a flattened interface for the AXI ports (see comments below).
  parameter type narrow_in_resp_flat_t = logic [$bits(narrow_in_resp_t)-1:0],
  parameter type narrow_out_req_flat_t = logic [$bits(narrow_out_req_t)-1:0],
  parameter type wide_out_req_flat_t   = logic [  $bits(wide_out_req_t)-1:0]
) (

  input  logic                                     soc_clk_i,
  input  logic                                     clu_clk_i,
  input  logic                                     rst_ni,
  input  logic                                     widemem_bypass_i,
  //-----------------------------
  // Interrupt ports
  //-----------------------------
  input  logic                 [      NrCores-1:0] debug_req_i,
  input  logic                 [      NrCores-1:0] meip_i,
  input  logic                 [      NrCores-1:0] mtip_i,
  input  logic                 [      NrCores-1:0] msip_i,
  //-----------------------------
  // Cluster base addressing
  //-----------------------------
  input  logic                 [              9:0] hart_base_id_i,
  input  logic                 [Cfg.AddrWidth-1:0] cluster_base_addr_i,
  input  logic                 [             31:0] boot_addr_i,
  //-----------------------------
  // Narrow AXI ports
  //-----------------------------
  input  narrow_in_req_t                           narrow_in_req_i,
  output narrow_in_resp_flat_t                     narrow_in_resp_flat_o,
  output narrow_out_req_flat_t [              1:0] narrow_out_req_flat_o,
  input  narrow_out_resp_t     [              1:0] narrow_out_resp_i,
  //-----------------------------
  //Wide AXI ports
  //-----------------------------
  output wide_out_req_flat_t                       wide_out_req_flat_o,
  input  wide_out_resp_t                           wide_out_resp_i
);

  `include "axi/typedef.svh"

  /* ------------------------------------------------------------------------------- */
  /*           Flattened interface signals for UPF structure workaround              */
  /* ------------------------------------------------------------------------------- */
  //
  // The UPF standard supported by QuestaSim cannot apply isolation strategies to
  // ports with "complex" types, such as AXI ports, which are structures.
  // To address this issue, at the interface of each power domain, signals are flattened
  // (e.g., narrow_in_resp_flat_o) and then internally reassigned to new structured signals
  // (e.g., narrow_in_resp_s), which can be propagated to downstream modules.
  //
  narrow_out_req_t [1:0] narrow_out_req_s;
  narrow_in_resp_t       narrow_in_resp_s;
  wide_out_req_t         wide_out_req_s;

  assign narrow_out_req_flat_o = narrow_out_req_s;
  assign narrow_in_resp_flat_o = narrow_in_resp_s;
  assign wide_out_req_flat_o   = wide_out_req_s;

  /* ------------------------------------------------------------------------------- */
  /* ------------------------------------------------------------------------------- */

  localparam int WideDataWidth = $bits(wide_out_req_s.w.data);

  localparam int WideMasterIdWidth = $bits(wide_out_req_s.aw.id);
  localparam int WideSlaveIdWidth = WideMasterIdWidth + $clog2(Cfg.AxiExtNumWideMst) - 1;

  localparam int NarrowSlaveIdWidth = $bits(narrow_in_req_i.aw.id);
  localparam int NarrowMasterIdWidth = $bits(narrow_out_req_s[0].aw.id);

  typedef logic [Cfg.AddrWidth-1:0] axi_addr_t;
  typedef logic [Cfg.AxiUserWidth-1:0] axi_user_t;

  typedef logic [Cfg.AxiDataWidth-1:0] axi_soc_data_narrow_t;
  typedef logic [Cfg.AxiDataWidth/8-1:0] axi_soc_strb_narrow_t;

  typedef logic [ClusterDataWidth-1:0] axi_cluster_data_narrow_t;
  typedef logic [ClusterDataWidth/8-1:0] axi_cluster_strb_narrow_t;

  typedef logic [WideDataWidth-1:0] axi_cluster_data_wide_t;
  typedef logic [WideDataWidth/8-1:0] axi_cluster_strb_wide_t;

  typedef logic [ClusterNarrowAxiMstIdWidth-1:0] axi_cluster_mst_id_width_narrow_t;
  typedef logic [ClusterNarrowAxiMstIdWidth-1+2:0] axi_cluster_slv_id_width_narrow_t;

  typedef logic [NarrowMasterIdWidth-1:0] axi_soc_mst_id_width_narrow_t;
  typedef logic [NarrowSlaveIdWidth-1:0] axi_soc_slv_id_width_narrow_t;

  typedef logic [WideMasterIdWidth-1:0] axi_mst_id_width_wide_t;
  typedef logic [WideMasterIdWidth-1+2:0] axi_slv_id_width_wide_t;

  `AXI_TYPEDEF_ALL(axi_cluster_out_wide, axi_addr_t, axi_slv_id_width_wide_t,
                   axi_cluster_data_wide_t, axi_cluster_strb_wide_t, axi_user_t)
  `AXI_TYPEDEF_ALL(axi_cluster_in_wide, axi_addr_t, axi_mst_id_width_wide_t,
                   axi_cluster_data_wide_t, axi_cluster_strb_wide_t, axi_user_t)

  `AXI_TYPEDEF_ALL(axi_soc_out_narrow, axi_addr_t, axi_soc_slv_id_width_narrow_t,
                   axi_soc_data_narrow_t, axi_soc_strb_narrow_t, axi_user_t)
  `AXI_TYPEDEF_ALL(axi_soc_in_narrow, axi_addr_t, axi_soc_mst_id_width_narrow_t,
                   axi_soc_data_narrow_t, axi_soc_strb_narrow_t, axi_user_t)

  `AXI_TYPEDEF_ALL(axi_cluster_out_narrow, axi_addr_t, axi_cluster_slv_id_width_narrow_t,
                   axi_cluster_data_narrow_t, axi_cluster_strb_narrow_t, axi_user_t)
  `AXI_TYPEDEF_ALL(axi_cluster_in_narrow, axi_addr_t, axi_cluster_mst_id_width_narrow_t,
                   axi_cluster_data_narrow_t, axi_cluster_strb_narrow_t, axi_user_t)

  `AXI_TYPEDEF_ALL(axi_cluster_out_narrow_socIW, axi_addr_t, axi_soc_mst_id_width_narrow_t,
                   axi_cluster_data_narrow_t, axi_cluster_strb_narrow_t, axi_user_t)
  `AXI_TYPEDEF_ALL(axi_cluster_in_narrow_socIW, axi_addr_t, axi_soc_slv_id_width_narrow_t,
                   axi_cluster_data_narrow_t, axi_cluster_strb_narrow_t, axi_user_t)

  // Cluster-side in- and out- narrow ports used in chimera adapter
  axi_cluster_in_narrow_req_t               clu_axi_adapter_slv_req;
  axi_cluster_in_narrow_resp_t              clu_axi_adapter_slv_resp;
  axi_cluster_out_narrow_req_t              clu_axi_adapter_mst_req;
  axi_cluster_out_narrow_resp_t             clu_axi_adapter_mst_resp;

  // Cluster-side in- and out- narrow ports used in narrow adapter
  axi_cluster_in_narrow_socIW_req_t         clu_axi_narrow_slv_req;
  axi_cluster_in_narrow_socIW_resp_t        clu_axi_narrow_slv_rsp;
  axi_cluster_out_narrow_socIW_req_t  [1:0] clu_axi_narrow_mst_req;
  axi_cluster_out_narrow_socIW_resp_t [1:0] clu_axi_narrow_mst_rsp;

  // Cluster-side out wide ports
  axi_cluster_out_wide_req_t                clu_axi_wide_mst_req;
  axi_cluster_out_wide_resp_t               clu_axi_wide_mst_resp;


  if (ClusterDataWidth != Cfg.AxiDataWidth) begin : gen_narrow_adapter

    narrow_adapter #(
      .narrow_in_req_t  (axi_soc_out_narrow_req_t),
      .narrow_in_resp_t (axi_soc_out_narrow_resp_t),
      .narrow_out_req_t (axi_soc_in_narrow_req_t),
      .narrow_out_resp_t(axi_soc_in_narrow_resp_t),

      .clu_narrow_in_req_t  (axi_cluster_in_narrow_socIW_req_t),
      .clu_narrow_in_resp_t (axi_cluster_in_narrow_socIW_resp_t),
      .clu_narrow_out_req_t (axi_cluster_out_narrow_socIW_req_t),
      .clu_narrow_out_resp_t(axi_cluster_out_narrow_socIW_resp_t),

      .MstPorts(2),
      .SlvPorts(1)

    ) i_cluster_narrow_adapter (
      .soc_clk_i(soc_clk_i),
      .rst_ni,

      // SoC side narrow.
      .narrow_in_req_i  (narrow_in_req_i),
      .narrow_in_resp_o (narrow_in_resp_s),
      .narrow_out_req_o (narrow_out_req_s),
      .narrow_out_resp_i(narrow_out_resp_i),

      // Cluster side narrow
      .clu_narrow_in_req_o  (clu_axi_narrow_slv_req),
      .clu_narrow_in_resp_i (clu_axi_narrow_slv_rsp),
      .clu_narrow_out_req_i (clu_axi_narrow_mst_req),
      .clu_narrow_out_resp_o(clu_axi_narrow_mst_rsp)

    );

  end else begin : gen_skip_narrow_adapter  // if (ClusterDataWidth != Cfg.AxiDataWidth)

    assign clu_axi_narrow_slv_req = narrow_in_req_i;
    assign narrow_in_resp_s       = clu_axi_narrow_slv_rsp;
    assign narrow_out_req_s       = clu_axi_narrow_mst_req;
    assign clu_axi_narrow_mst_rsp = narrow_out_resp_i;

  end

  chimera_cluster_adapter #(
    .WidePassThroughRegionStart(Cfg.MemIslRegionStart),
    .WidePassThroughRegionEnd  (Cfg.MemIslRegionEnd),

    .narrow_in_req_t  (axi_cluster_in_narrow_socIW_req_t),
    .narrow_in_resp_t (axi_cluster_in_narrow_socIW_resp_t),
    .narrow_out_req_t (axi_cluster_out_narrow_socIW_req_t),
    .narrow_out_resp_t(axi_cluster_out_narrow_socIW_resp_t),

    .clu_narrow_in_req_t  (axi_cluster_in_narrow_req_t),
    .clu_narrow_in_resp_t (axi_cluster_in_narrow_resp_t),
    .clu_narrow_out_req_t (axi_cluster_out_narrow_req_t),
    .clu_narrow_out_resp_t(axi_cluster_out_narrow_resp_t),

    .wide_out_req_t (wide_out_req_t),
    .wide_out_resp_t(wide_out_resp_t),

    .clu_wide_out_req_t (axi_cluster_out_wide_req_t),
    .clu_wide_out_resp_t(axi_cluster_out_wide_resp_t)

  ) i_cluster_axi_adapter (
    .soc_clk_i(soc_clk_i),
    .clu_clk_i(clu_clk_i),
    .rst_ni,

    .narrow_in_req_i  (clu_axi_narrow_slv_req),
    .narrow_in_resp_o (clu_axi_narrow_slv_rsp),
    .narrow_out_req_o (clu_axi_narrow_mst_req),
    .narrow_out_resp_i(clu_axi_narrow_mst_rsp),

    .clu_narrow_in_req_o  (clu_axi_adapter_slv_req),
    .clu_narrow_in_resp_i (clu_axi_adapter_slv_resp),
    .clu_narrow_out_req_i (clu_axi_adapter_mst_req),
    .clu_narrow_out_resp_o(clu_axi_adapter_mst_resp),

    .wide_out_req_o     (wide_out_req_s),
    .wide_out_resp_i    (wide_out_resp_i),
    .clu_wide_out_req_i (clu_axi_wide_mst_req),
    .clu_wide_out_resp_o(clu_axi_wide_mst_resp),

    .wide_mem_bypass_mode_i(widemem_bypass_i)
  );

  typedef struct packed {
    logic [2:0] ema;
    logic [1:0] emaw;
    logic [0:0] emas;
  } sram_cfg_t;

  typedef struct packed {
    sram_cfg_t icache_tag;
    sram_cfg_t icache_data;
    sram_cfg_t tcdm;
  } sram_cfgs_t;

  localparam int unsigned NumIntOutstandingLoads[NrCores] = '{NrCores{32'h1}};
  localparam int unsigned NumIntOutstandingMem[NrCores] = '{NrCores{32'h4}};

  snitch_cluster #(
    .PhysicalAddrWidth(Cfg.AddrWidth),
    .NarrowDataWidth  (ClusterDataWidth),            // SCHEREMO: Convolve needs this...
    .WideDataWidth    (WideDataWidth),
    .NarrowIdWidthIn  (ClusterNarrowAxiMstIdWidth),
    .WideIdWidthIn    (WideMasterIdWidth),
    .NarrowUserWidth  (Cfg.AxiUserWidth),
    .WideUserWidth    (Cfg.AxiUserWidth),

    .BootAddr(SnitchBootROMRegionStart),

    .NrHives          (1),
    .NrCores          (NrCores),
    .TCDMDepth        (1024),
    .ZeroMemorySize   (64),
    .ClusterPeriphSize(64),
    .NrBanks          (16),

    .DMANumAxInFlight(3),
    .DMAReqFifoDepth (3),

    .ICacheLineWidth('{256}),
    .ICacheLineCount('{16}),
    .ICacheSets     ('{2}),

    .VMSupport(0),
    .Xdma     ({1'b1, {(NrCores - 1) {1'b0}}}),

    .NumIntOutstandingLoads(NumIntOutstandingLoads),
    .NumIntOutstandingMem  (NumIntOutstandingMem),
    .RegisterOffloadReq    (1),
    .RegisterOffloadRsp    (1),
    .RegisterCoreReq       (1),
    .RegisterCoreRsp       (1),

    .narrow_in_req_t (axi_cluster_in_narrow_req_t),
    .narrow_in_resp_t(axi_cluster_in_narrow_resp_t),
    .wide_in_req_t   (axi_cluster_in_wide_req_t),
    .wide_in_resp_t  (axi_cluster_in_wide_resp_t),

    .narrow_out_req_t (axi_cluster_out_narrow_req_t),
    .narrow_out_resp_t(axi_cluster_out_narrow_resp_t),
    .wide_out_req_t   (axi_cluster_out_wide_req_t),
    .wide_out_resp_t  (axi_cluster_out_wide_resp_t),

    .sram_cfg_t (sram_cfg_t),
    .sram_cfgs_t(sram_cfgs_t),

    .RegisterExtWide  ('0),
    .RegisterExtNarrow('0)
  ) i_test_cluster (

    .clk_i          (clu_clk_i),
    .clk_d2_bypass_i('0),
    .rst_ni,

    .debug_req_i(debug_req_i),
    .meip_i     (meip_i),
    .mtip_i     (mtip_i),
    .msip_i     (msip_i),

    .hart_base_id_i     (hart_base_id_i),
    .cluster_base_addr_i(cluster_base_addr_i),
    .sram_cfgs_i        ('0),

    .narrow_in_req_i  (clu_axi_adapter_slv_req),
    .narrow_in_resp_o (clu_axi_adapter_slv_resp),
    .narrow_out_req_o (clu_axi_adapter_mst_req),
    .narrow_out_resp_i(clu_axi_adapter_mst_resp),
    .wide_in_req_i    ('0),
    .wide_in_resp_o   (),
    .wide_out_req_o   (clu_axi_wide_mst_req),
    .wide_out_resp_i  (clu_axi_wide_mst_resp)

  );
endmodule

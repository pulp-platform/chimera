// Copyright 2022 ETH Zurich and University of Bologna.
// Solderpad Hardware License, Version 0.51, see LICENSE for details.
// SPDX-License-Identifier: SHL-0.51
//
// Fabian Schuiki <fschuiki@iis.ee.ethz.ch>
// Florian Zaruba <zarubaf@iis.ee.ethz.ch>
// Stefan Mach <smach@iis.ee.ethz.ch>
// Thomas Benz <tbenz@iis.ee.ethz.ch>
// Paul Scheffler <paulsc@iis.ee.ethz.ch>
// Wolfgang Roenninger <wroennin@iis.ee.ethz.ch>
//
// AUTOMATICALLY GENERATED by gen_bootrom.py; edit the script instead.

module snitch_bootrom #(
    parameter int unsigned AddrWidth = 32,
    parameter int unsigned DataWidth = 32
)(
    input  logic                 clk_i,
    input  logic                 rst_ni,
    input  logic                 req_i,
    input  logic [AddrWidth-1:0] addr_i,
    output logic [DataWidth-1:0] data_o
);
    localparam unsigned NumWords = 128;
    logic [$clog2(NumWords)-1:0] word;

    assign word = addr_i / (DataWidth / 8);

    always_comb begin
        data_o = '0;
        unique case (word)
        000: data_o = 32'h30057073 /* 0x0000 */;
            001: data_o = 32'h138000ef /* 0x0004 */;
            002: data_o = 32'h00000297 /* 0x0008 */;
            003: data_o = 32'h09828293 /* 0x000c */;
            004: data_o = 32'h30529073 /* 0x0010 */;
            005: data_o = 32'h00000293 /* 0x0014 */;
            006: data_o = 32'h00000313 /* 0x0018 */;
            007: data_o = 32'h00000393 /* 0x001c */;
            008: data_o = 32'h00000413 /* 0x0020 */;
            009: data_o = 32'h00000493 /* 0x0024 */;
            010: data_o = 32'h00000513 /* 0x0028 */;
            011: data_o = 32'h00000593 /* 0x002c */;
            012: data_o = 32'h00000613 /* 0x0030 */;
            013: data_o = 32'h00000693 /* 0x0034 */;
            014: data_o = 32'h00000713 /* 0x0038 */;
            015: data_o = 32'h00000793 /* 0x003c */;
            016: data_o = 32'h00000813 /* 0x0040 */;
            017: data_o = 32'h00000893 /* 0x0044 */;
            018: data_o = 32'h00000913 /* 0x0048 */;
            019: data_o = 32'h00000993 /* 0x004c */;
            020: data_o = 32'h00000a13 /* 0x0050 */;
            021: data_o = 32'h00000a93 /* 0x0054 */;
            022: data_o = 32'h00000b13 /* 0x0058 */;
            023: data_o = 32'h00000b93 /* 0x005c */;
            024: data_o = 32'h00000c13 /* 0x0060 */;
            025: data_o = 32'h00000c93 /* 0x0064 */;
            026: data_o = 32'h00000d13 /* 0x0068 */;
            027: data_o = 32'h00000d93 /* 0x006c */;
            028: data_o = 32'h00000e13 /* 0x0070 */;
            029: data_o = 32'h00000e93 /* 0x0074 */;
            030: data_o = 32'h00000f13 /* 0x0078 */;
            031: data_o = 32'h00000f93 /* 0x007c */;
            032: data_o = 32'h10500073 /* 0x0080 */;
            033: data_o = 32'h00001297 /* 0x0084 */;
            034: data_o = 32'hf7c28293 /* 0x0088 */;
            035: data_o = 32'h0002a283 /* 0x008c */;
            036: data_o = 32'h000280e7 /* 0x0090 */;
            037: data_o = 32'h02c000ef /* 0x0094 */;
            038: data_o = 32'hf7dff06f /* 0x0098 */;
            039: data_o = 32'h00000013 /* 0x009c */;
            040: data_o = 32'h00001297 /* 0x00a0 */;
            041: data_o = 32'hf6028293 /* 0x00a4 */;
            042: data_o = 32'h0042a283 /* 0x00a8 */;
            043: data_o = 32'h000280e7 /* 0x00ac */;
            044: data_o = 32'h30200073 /* 0x00b0 */;
            045: data_o = 32'h00000000 /* 0x00b4 */;
            046: data_o = 32'h00000000 /* 0x00b8 */;
            047: data_o = 32'h00000000 /* 0x00bc */;
            048: data_o = 32'hf14027f3 /* 0x00c0 */;
            049: data_o = 32'h01300713 /* 0x00c4 */;
            050: data_o = 32'h0ff7f793 /* 0x00c8 */;
            051: data_o = 32'h00156513 /* 0x00cc */;
            052: data_o = 32'h04e78463 /* 0x00d0 */;
            053: data_o = 32'h00f76c63 /* 0x00d4 */;
            054: data_o = 32'h00100713 /* 0x00d8 */;
            055: data_o = 32'h02e78263 /* 0x00dc */;
            056: data_o = 32'h00a00713 /* 0x00e0 */;
            057: data_o = 32'h02e78463 /* 0x00e4 */;
            058: data_o = 32'h00008067 /* 0x00e8 */;
            059: data_o = 32'h01c00713 /* 0x00ec */;
            060: data_o = 32'h02e78a63 /* 0x00f0 */;
            061: data_o = 32'h02500713 /* 0x00f4 */;
            062: data_o = 32'h02e78c63 /* 0x00f8 */;
            063: data_o = 32'h00008067 /* 0x00fc */;
            064: data_o = 32'h300017b7 /* 0x0100 */;
            065: data_o = 32'h00a7a423 /* 0x0104 */;
            066: data_o = 32'h00008067 /* 0x0108 */;
            067: data_o = 32'h300017b7 /* 0x010c */;
            068: data_o = 32'h00a7a623 /* 0x0110 */;
            069: data_o = 32'h00008067 /* 0x0114 */;
            070: data_o = 32'h300017b7 /* 0x0118 */;
            071: data_o = 32'h00a7a823 /* 0x011c */;
            072: data_o = 32'h00008067 /* 0x0120 */;
            073: data_o = 32'h300017b7 /* 0x0124 */;
            074: data_o = 32'h00a7aa23 /* 0x0128 */;
            075: data_o = 32'h00008067 /* 0x012c */;
            076: data_o = 32'h300017b7 /* 0x0130 */;
            077: data_o = 32'h00a7ac23 /* 0x0134 */;
            078: data_o = 32'h00008067 /* 0x0138 */;
            079: data_o = 32'h304467f3 /* 0x013c */;
            080: data_o = 32'h300467f3 /* 0x0140 */;
            081: data_o = 32'h00008067 /* 0x0144 */;
            082: data_o = 32'h00000000 /* 0x0148 */;
            083: data_o = 32'h00000000 /* 0x014c */;
            084: data_o = 32'h00000000 /* 0x0150 */;
            085: data_o = 32'h00000000 /* 0x0154 */;
            086: data_o = 32'h00000000 /* 0x0158 */;
            087: data_o = 32'h00000000 /* 0x015c */;
            088: data_o = 32'h00000000 /* 0x0160 */;
            089: data_o = 32'h00000000 /* 0x0164 */;
            090: data_o = 32'h00000000 /* 0x0168 */;
            091: data_o = 32'h00000000 /* 0x016c */;
            092: data_o = 32'h00000000 /* 0x0170 */;
            093: data_o = 32'h00000000 /* 0x0174 */;
            094: data_o = 32'h00000000 /* 0x0178 */;
            095: data_o = 32'h00000000 /* 0x017c */;
            096: data_o = 32'h00000000 /* 0x0180 */;
            097: data_o = 32'h00000000 /* 0x0184 */;
            098: data_o = 32'h00000000 /* 0x0188 */;
            099: data_o = 32'h00000000 /* 0x018c */;
            100: data_o = 32'h00000000 /* 0x0190 */;
            101: data_o = 32'h00000000 /* 0x0194 */;
            102: data_o = 32'h00000000 /* 0x0198 */;
            103: data_o = 32'h00000000 /* 0x019c */;
            104: data_o = 32'h00000000 /* 0x01a0 */;
            105: data_o = 32'h00000000 /* 0x01a4 */;
            106: data_o = 32'h00000000 /* 0x01a8 */;
            107: data_o = 32'h00000000 /* 0x01ac */;
            108: data_o = 32'h00000000 /* 0x01b0 */;
            109: data_o = 32'h00000000 /* 0x01b4 */;
            110: data_o = 32'h00000000 /* 0x01b8 */;
            111: data_o = 32'h00000000 /* 0x01bc */;
            112: data_o = 32'h00000000 /* 0x01c0 */;
            113: data_o = 32'h00000000 /* 0x01c4 */;
            114: data_o = 32'h00000000 /* 0x01c8 */;
            115: data_o = 32'h00000000 /* 0x01cc */;
            116: data_o = 32'h00000000 /* 0x01d0 */;
            117: data_o = 32'h00000000 /* 0x01d4 */;
            118: data_o = 32'h00000000 /* 0x01d8 */;
            119: data_o = 32'h00000000 /* 0x01dc */;
            120: data_o = 32'h00000000 /* 0x01e0 */;
            121: data_o = 32'h00000000 /* 0x01e4 */;
            122: data_o = 32'h00000000 /* 0x01e8 */;
            123: data_o = 32'h00000000 /* 0x01ec */;
            124: data_o = 32'h00000000 /* 0x01f0 */;
            125: data_o = 32'h00000000 /* 0x01f4 */;
            126: data_o = 32'h00000000 /* 0x01f8 */;
            127: data_o = 32'h00000000 /* 0x01fc */;
            default: data_o = '0;
        endcase
    end

endmodule

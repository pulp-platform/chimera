// Copyright 2023 ETH Zurich and University of Bologna.
// Solderpad Hardware License, Version 0.51, see LICENSE for details.
// SPDX-License-Identifier: SHL-0.51
//
// Yvan Tortorella <yvan.tortorella@unibo.it>

`include "register_interface/typedef.svh"

module hyperbus_wrap #(
  parameter int unsigned NumChips = -1,
  parameter int unsigned NumPhys = 2,
  parameter int unsigned IsClockODelayed = 0,
  parameter int unsigned AxiAddrWidth = -1,
  parameter int unsigned AxiDataWidth = -1,
  parameter int unsigned AxiIdWidth = -1,
  parameter int unsigned AxiUserWidth = -1,
  parameter int unsigned AxiMaxTrans = 0,
  parameter type axi_req_t = logic,
  parameter type axi_rsp_t = logic,
  parameter type axi_w_chan_t = logic,
  parameter type axi_b_chan_t = logic,
  parameter type axi_ar_chan_t = logic,
  parameter type axi_r_chan_t = logic,
  parameter type axi_aw_chan_t = logic,
  parameter int unsigned RegAddrWidth = -1,
  parameter int unsigned RegDataWidth = -1,
  parameter type reg_req_t = logic,
  parameter type reg_rsp_t = logic,
  parameter type reg_addr_t = logic [RegAddrWidth-1:0],
  parameter type reg_data_t = logic [RegDataWidth-1:0],
  parameter type reg_strb_t = logic [RegDataWidth/8-1:0],
  // The below have sensible defaults, but should be set on integration!
  parameter int unsigned RxFifoLogDepth = 2,
  parameter int unsigned TxFifoLogDepth = 2,
  parameter logic [RegDataWidth-1:0] RstChipBase = 'h0,  // Base address for all chips
  parameter logic [RegDataWidth-1:0] RstChipSpace = 'h1_0000,  // 64 KiB: Current maximum H
                                                               // yperBus device size
  parameter int unsigned PhyStartupCycles = 300 * 200,  /* us*MHz */
  // Conservative maximum
  // frequency estimate
  parameter int unsigned AxiLogDepth = 3,
  parameter int unsigned AxiSlaveArWidth = 0,
  parameter int unsigned AxiSlaveAwWidth = 0,
  parameter int unsigned AxiSlaveBWidth = 0,
  parameter int unsigned AxiSlaveRWidth = 0,
  parameter int unsigned AxiSlaveWWidth = 0,
  parameter int unsigned CdcSyncStages = 0
) (
  input  logic                                          clk_i,
  input  logic                                          rst_ni,
  input  logic                                          test_mode_i,
  // AXI bus
  input  logic      [AxiSlaveArWidth-1:0]               axi_slave_ar_data_i,
  input  logic      [      AxiLogDepth:0]               axi_slave_ar_wptr_i,
  output logic      [      AxiLogDepth:0]               axi_slave_ar_rptr_o,
  input  logic      [AxiSlaveAwWidth-1:0]               axi_slave_aw_data_i,
  input  logic      [      AxiLogDepth:0]               axi_slave_aw_wptr_i,
  output logic      [      AxiLogDepth:0]               axi_slave_aw_rptr_o,
  output logic      [ AxiSlaveBWidth-1:0]               axi_slave_b_data_o,
  output logic      [      AxiLogDepth:0]               axi_slave_b_wptr_o,
  input  logic      [      AxiLogDepth:0]               axi_slave_b_rptr_i,
  output logic      [ AxiSlaveRWidth-1:0]               axi_slave_r_data_o,
  output logic      [      AxiLogDepth:0]               axi_slave_r_wptr_o,
  input  logic      [      AxiLogDepth:0]               axi_slave_r_rptr_i,
  input  logic      [ AxiSlaveWWidth-1:0]               axi_slave_w_data_i,
  input  logic      [      AxiLogDepth:0]               axi_slave_w_wptr_i,
  output logic      [      AxiLogDepth:0]               axi_slave_w_rptr_o,
  // Reg bus
  input  reg_addr_t                                     rbus_req_addr_i,
  input  logic                                          rbus_req_write_i,
  input  reg_data_t                                     rbus_req_wdata_i,
  input  reg_strb_t                                     rbus_req_wstrb_i,
  input  logic                                          rbus_req_valid_i,
  output reg_data_t                                     rbus_rsp_rdata_o,
  output logic                                          rbus_rsp_ready_o,
  output logic                                          rbus_rsp_error_o,
  // Physical interace: HyperBus PADs
  output logic      [        NumPhys-1:0][NumChips-1:0] hyper_cs_no,
  output logic      [        NumPhys-1:0]               hyper_ck_o,
  output logic      [        NumPhys-1:0]               hyper_ck_no,
  output logic      [        NumPhys-1:0]               hyper_rwds_o,
  input  logic      [        NumPhys-1:0]               hyper_rwds_i,
  output logic      [        NumPhys-1:0]               hyper_rwds_oe_o,
  input  logic      [        NumPhys-1:0][         7:0] hyper_dq_i,
  output logic      [        NumPhys-1:0][         7:0] hyper_dq_o,
  output logic      [        NumPhys-1:0]               hyper_dq_oe_o,
  output logic      [        NumPhys-1:0]               hyper_reset_no
);

  reg_req_t reg_req;
  reg_rsp_t reg_rsp;

  typedef struct packed {
    logic [31:0]             idx;
    logic [AxiAddrWidth-1:0] start_addr;
    logic [AxiAddrWidth-1:0] end_addr;
  } addr_rule_t;

  axi_req_t hyper_req;
  axi_rsp_t hyper_rsp;

  axi_cdc_dst #(
    .LogDepth  (AxiLogDepth),
    .SyncStages(CdcSyncStages),
    .aw_chan_t (axi_aw_chan_t),
    .w_chan_t  (axi_w_chan_t),
    .b_chan_t  (axi_b_chan_t),
    .ar_chan_t (axi_ar_chan_t),
    .r_chan_t  (axi_r_chan_t),
    .axi_req_t (axi_req_t),
    .axi_resp_t(axi_rsp_t)
  ) i_hyper_cdc_dst (
    // asynchronous slave port
    .async_data_slave_aw_data_i(axi_slave_aw_data_i),
    .async_data_slave_aw_wptr_i(axi_slave_aw_wptr_i),
    .async_data_slave_aw_rptr_o(axi_slave_aw_rptr_o),
    .async_data_slave_w_data_i (axi_slave_w_data_i),
    .async_data_slave_w_wptr_i (axi_slave_w_wptr_i),
    .async_data_slave_w_rptr_o (axi_slave_w_rptr_o),
    .async_data_slave_b_data_o (axi_slave_b_data_o),
    .async_data_slave_b_wptr_o (axi_slave_b_wptr_o),
    .async_data_slave_b_rptr_i (axi_slave_b_rptr_i),
    .async_data_slave_ar_data_i(axi_slave_ar_data_i),
    .async_data_slave_ar_wptr_i(axi_slave_ar_wptr_i),
    .async_data_slave_ar_rptr_o(axi_slave_ar_rptr_o),
    .async_data_slave_r_data_o (axi_slave_r_data_o),
    .async_data_slave_r_wptr_o (axi_slave_r_wptr_o),
    .async_data_slave_r_rptr_i (axi_slave_r_rptr_i),
    // synchronous master port
    .dst_clk_i                 (clk_i),
    .dst_rst_ni                (rst_ni),
    .dst_req_o                 (hyper_req),
    .dst_resp_i                (hyper_rsp)
  );

  assign reg_req.addr     = rbus_req_addr_i;
  assign reg_req.write    = rbus_req_write_i;
  assign reg_req.wdata    = rbus_req_wdata_i;
  assign reg_req.wstrb    = rbus_req_wstrb_i;
  assign reg_req.valid    = rbus_req_valid_i;
  assign rbus_rsp_rdata_o = reg_rsp.rdata;
  assign rbus_rsp_ready_o = reg_rsp.ready;
  assign rbus_rsp_error_o = reg_rsp.error;

  hyperbus #(
    .NumChips        (NumChips),
    .NumPhys         (NumPhys),
    .IsClockODelayed (IsClockODelayed),
    .AxiAddrWidth    (AxiAddrWidth),
    .AxiDataWidth    (AxiDataWidth),
    .AxiIdWidth      (AxiIdWidth),
    .AxiUserWidth    (AxiUserWidth),
    .axi_req_t       (axi_req_t),
    .axi_rsp_t       (axi_rsp_t),
    .RegAddrWidth    (RegAddrWidth),
    .RegDataWidth    (RegDataWidth),
    .reg_req_t       (reg_req_t),
    .reg_rsp_t       (reg_rsp_t),
    .axi_rule_t      (addr_rule_t),
    .RxFifoLogDepth  (RxFifoLogDepth),
    .TxFifoLogDepth  (TxFifoLogDepth),
    .RstChipBase     (RstChipBase),
    .RstChipSpace    (RstChipSpace),
    .PhyStartupCycles(PhyStartupCycles),
    .AxiLogDepth     (AxiLogDepth),
    .SyncStages      (CdcSyncStages)
  ) i_hyperbus (
    .clk_phy_i  (clk_i),
    .rst_phy_ni (rst_ni),
    .clk_sys_i  (clk_i),
    .rst_sys_ni (rst_ni),
    .test_mode_i(test_mode_i),
    .axi_req_i  (hyper_req),
    .axi_rsp_o  (hyper_rsp),
    .reg_req_i  (reg_req),
    .reg_rsp_o  (reg_rsp),
    .hyper_cs_no,
    .hyper_ck_o,
    .hyper_ck_no,
    .hyper_rwds_o,
    .hyper_rwds_i,
    .hyper_rwds_oe_o,
    .hyper_dq_i,
    .hyper_dq_o,
    .hyper_dq_oe_o,
    .hyper_reset_no
  );

endmodule : hyperbus_wrap

// Copyright 2022 ETH Zurich and University of Bologna.
// Solderpad Hardware License, Version 0.51, see LICENSE for details.
// SPDX-License-Identifier: SHL-0.51
//
// Fabian Schuiki <fschuiki@iis.ee.ethz.ch>
// Florian Zaruba <zarubaf@iis.ee.ethz.ch>
// Stefan Mach <smach@iis.ee.ethz.ch>
// Thomas Benz <tbenz@iis.ee.ethz.ch>
// Paul Scheffler <paulsc@iis.ee.ethz.ch>
// Wolfgang Roenninger <wroennin@iis.ee.ethz.ch>
//
// AUTOMATICALLY GENERATED by gen_bootrom.py; edit the script instead.

module snitch_bootrom #(
    parameter int unsigned AddrWidth = 32,
    parameter int unsigned DataWidth = 32
)(
    input  logic                 clk_i,
    input  logic                 rst_ni,
    input  logic                 req_i,
    input  logic [AddrWidth-1:0] addr_i,
    output logic [DataWidth-1:0] data_o
);
    localparam unsigned NumWords = 256;
    logic [$clog2(NumWords)-1:0] word;

    assign word = addr_i / (DataWidth / 8);

    always_comb begin
        data_o = '0;
        unique case (word)
        000: data_o = 32'h30057073 /* 0x0000 */;
            001: data_o = 32'h00000097 /* 0x0004 */;
            002: data_o = 32'h22c080e7 /* 0x0008 */;
            003: data_o = 32'h00000297 /* 0x000c */;
            004: data_o = 32'h0b428293 /* 0x0010 */;
            005: data_o = 32'h30529073 /* 0x0014 */;
            006: data_o = 32'h00000293 /* 0x0018 */;
            007: data_o = 32'h00000313 /* 0x001c */;
            008: data_o = 32'h00000393 /* 0x0020 */;
            009: data_o = 32'h00000413 /* 0x0024 */;
            010: data_o = 32'h00000493 /* 0x0028 */;
            011: data_o = 32'h00000513 /* 0x002c */;
            012: data_o = 32'h00000593 /* 0x0030 */;
            013: data_o = 32'h00000613 /* 0x0034 */;
            014: data_o = 32'h00000693 /* 0x0038 */;
            015: data_o = 32'h00000713 /* 0x003c */;
            016: data_o = 32'h00000793 /* 0x0040 */;
            017: data_o = 32'h00000813 /* 0x0044 */;
            018: data_o = 32'h00000893 /* 0x0048 */;
            019: data_o = 32'h00000913 /* 0x004c */;
            020: data_o = 32'h00000993 /* 0x0050 */;
            021: data_o = 32'h00000a13 /* 0x0054 */;
            022: data_o = 32'h00000a93 /* 0x0058 */;
            023: data_o = 32'h00000b13 /* 0x005c */;
            024: data_o = 32'h00000b93 /* 0x0060 */;
            025: data_o = 32'h00000c13 /* 0x0064 */;
            026: data_o = 32'h00000c93 /* 0x0068 */;
            027: data_o = 32'h00000d13 /* 0x006c */;
            028: data_o = 32'h00000d93 /* 0x0070 */;
            029: data_o = 32'h00000e13 /* 0x0074 */;
            030: data_o = 32'h00000e93 /* 0x0078 */;
            031: data_o = 32'h00000f13 /* 0x007c */;
            032: data_o = 32'h00000f93 /* 0x0080 */;
            033: data_o = 32'h00000097 /* 0x0084 */;
            034: data_o = 32'h0d8080e7 /* 0x0088 */;
            035: data_o = 32'h10500073 /* 0x008c */;
            036: data_o = 32'h00000097 /* 0x0090 */;
            037: data_o = 32'h050080e7 /* 0x0094 */;
            038: data_o = 32'h00001297 /* 0x0098 */;
            039: data_o = 32'hf6828293 /* 0x009c */;
            040: data_o = 32'h0002a283 /* 0x00a0 */;
            041: data_o = 32'h000280e7 /* 0x00a4 */;
            042: data_o = 32'h00000097 /* 0x00a8 */;
            043: data_o = 32'h11c080e7 /* 0x00ac */;
            044: data_o = 32'hf69ff06f /* 0x00b0 */;
            045: data_o = 32'h00000013 /* 0x00b4 */;
            046: data_o = 32'h00000013 /* 0x00b8 */;
            047: data_o = 32'h00000013 /* 0x00bc */;
            048: data_o = 32'h00001297 /* 0x00c0 */;
            049: data_o = 32'hf4028293 /* 0x00c4 */;
            050: data_o = 32'h0042a283 /* 0x00c8 */;
            051: data_o = 32'h000280e7 /* 0x00cc */;
            052: data_o = 32'h30200073 /* 0x00d0 */;
            053: data_o = 32'h00000000 /* 0x00d4 */;
            054: data_o = 32'h00000000 /* 0x00d8 */;
            055: data_o = 32'h00000000 /* 0x00dc */;
            056: data_o = 32'hf14027f3 /* 0x00e0 */;
            057: data_o = 32'hfff78793 /* 0x00e4 */;
            058: data_o = 32'h0ff7f793 /* 0x00e8 */;
            059: data_o = 32'h00800713 /* 0x00ec */;
            060: data_o = 32'h06f76463 /* 0x00f0 */;
            061: data_o = 32'h30000737 /* 0x00f4 */;
            062: data_o = 32'h00279793 /* 0x00f8 */;
            063: data_o = 32'h23c70713 /* 0x00fc */;
            064: data_o = 32'h00e787b3 /* 0x0100 */;
            065: data_o = 32'h0007a783 /* 0x0104 */;
            066: data_o = 32'h00078067 /* 0x0108 */;
            067: data_o = 32'h300017b7 /* 0x010c */;
            068: data_o = 32'h00100713 /* 0x0110 */;
            069: data_o = 32'h04e7a223 /* 0x0114 */;
            070: data_o = 32'h00008067 /* 0x0118 */;
            071: data_o = 32'h300017b7 /* 0x011c */;
            072: data_o = 32'h00100713 /* 0x0120 */;
            073: data_o = 32'h04e7a423 /* 0x0124 */;
            074: data_o = 32'h00008067 /* 0x0128 */;
            075: data_o = 32'h300017b7 /* 0x012c */;
            076: data_o = 32'h00100713 /* 0x0130 */;
            077: data_o = 32'h04e7a623 /* 0x0134 */;
            078: data_o = 32'h00008067 /* 0x0138 */;
            079: data_o = 32'h300017b7 /* 0x013c */;
            080: data_o = 32'h00100713 /* 0x0140 */;
            081: data_o = 32'h04e7a823 /* 0x0144 */;
            082: data_o = 32'h00008067 /* 0x0148 */;
            083: data_o = 32'h300017b7 /* 0x014c */;
            084: data_o = 32'h00100713 /* 0x0150 */;
            085: data_o = 32'h04e7aa23 /* 0x0154 */;
            086: data_o = 32'h00008067 /* 0x0158 */;
            087: data_o = 32'hf14027f3 /* 0x015c */;
            088: data_o = 32'hfff78793 /* 0x0160 */;
            089: data_o = 32'h0ff7f793 /* 0x0164 */;
            090: data_o = 32'h00800713 /* 0x0168 */;
            091: data_o = 32'h04f76a63 /* 0x016c */;
            092: data_o = 32'h30000737 /* 0x0170 */;
            093: data_o = 32'h00279793 /* 0x0174 */;
            094: data_o = 32'h26070713 /* 0x0178 */;
            095: data_o = 32'h00e787b3 /* 0x017c */;
            096: data_o = 32'h0007a783 /* 0x0180 */;
            097: data_o = 32'h00078067 /* 0x0184 */;
            098: data_o = 32'h300017b7 /* 0x0188 */;
            099: data_o = 32'h0407a223 /* 0x018c */;
            100: data_o = 32'h00008067 /* 0x0190 */;
            101: data_o = 32'h300017b7 /* 0x0194 */;
            102: data_o = 32'h0407a423 /* 0x0198 */;
            103: data_o = 32'h00008067 /* 0x019c */;
            104: data_o = 32'h300017b7 /* 0x01a0 */;
            105: data_o = 32'h0407a623 /* 0x01a4 */;
            106: data_o = 32'h00008067 /* 0x01a8 */;
            107: data_o = 32'h300017b7 /* 0x01ac */;
            108: data_o = 32'h0407a823 /* 0x01b0 */;
            109: data_o = 32'h00008067 /* 0x01b4 */;
            110: data_o = 32'h300017b7 /* 0x01b8 */;
            111: data_o = 32'h0407aa23 /* 0x01bc */;
            112: data_o = 32'h00008067 /* 0x01c0 */;
            113: data_o = 32'hf14027f3 /* 0x01c4 */;
            114: data_o = 32'hfff78793 /* 0x01c8 */;
            115: data_o = 32'h0ff7f793 /* 0x01cc */;
            116: data_o = 32'h00800713 /* 0x01d0 */;
            117: data_o = 32'h00156513 /* 0x01d4 */;
            118: data_o = 32'h04f76a63 /* 0x01d8 */;
            119: data_o = 32'h30000737 /* 0x01dc */;
            120: data_o = 32'h00279793 /* 0x01e0 */;
            121: data_o = 32'h28470713 /* 0x01e4 */;
            122: data_o = 32'h00e787b3 /* 0x01e8 */;
            123: data_o = 32'h0007a783 /* 0x01ec */;
            124: data_o = 32'h00078067 /* 0x01f0 */;
            125: data_o = 32'h300017b7 /* 0x01f4 */;
            126: data_o = 32'h00a7a423 /* 0x01f8 */;
            127: data_o = 32'h00008067 /* 0x01fc */;
            128: data_o = 32'h300017b7 /* 0x0200 */;
            129: data_o = 32'h00a7a623 /* 0x0204 */;
            130: data_o = 32'h00008067 /* 0x0208 */;
            131: data_o = 32'h300017b7 /* 0x020c */;
            132: data_o = 32'h00a7a823 /* 0x0210 */;
            133: data_o = 32'h00008067 /* 0x0214 */;
            134: data_o = 32'h300017b7 /* 0x0218 */;
            135: data_o = 32'h00a7aa23 /* 0x021c */;
            136: data_o = 32'h00008067 /* 0x0220 */;
            137: data_o = 32'h300017b7 /* 0x0224 */;
            138: data_o = 32'h00a7ac23 /* 0x0228 */;
            139: data_o = 32'h00008067 /* 0x022c */;
            140: data_o = 32'h304467f3 /* 0x0230 */;
            141: data_o = 32'h300467f3 /* 0x0234 */;
            142: data_o = 32'h00008067 /* 0x0238 */;
            143: data_o = 32'h3000010c /* 0x023c */;
            144: data_o = 32'h30000158 /* 0x0240 */;
            145: data_o = 32'h3000011c /* 0x0244 */;
            146: data_o = 32'h30000158 /* 0x0248 */;
            147: data_o = 32'h3000012c /* 0x024c */;
            148: data_o = 32'h30000158 /* 0x0250 */;
            149: data_o = 32'h3000013c /* 0x0254 */;
            150: data_o = 32'h30000158 /* 0x0258 */;
            151: data_o = 32'h3000014c /* 0x025c */;
            152: data_o = 32'h30000188 /* 0x0260 */;
            153: data_o = 32'h300001c0 /* 0x0264 */;
            154: data_o = 32'h30000194 /* 0x0268 */;
            155: data_o = 32'h300001c0 /* 0x026c */;
            156: data_o = 32'h300001a0 /* 0x0270 */;
            157: data_o = 32'h300001c0 /* 0x0274 */;
            158: data_o = 32'h300001ac /* 0x0278 */;
            159: data_o = 32'h300001c0 /* 0x027c */;
            160: data_o = 32'h300001b8 /* 0x0280 */;
            161: data_o = 32'h300001f4 /* 0x0284 */;
            162: data_o = 32'h3000022c /* 0x0288 */;
            163: data_o = 32'h30000200 /* 0x028c */;
            164: data_o = 32'h3000022c /* 0x0290 */;
            165: data_o = 32'h3000020c /* 0x0294 */;
            166: data_o = 32'h3000022c /* 0x0298 */;
            167: data_o = 32'h30000218 /* 0x029c */;
            168: data_o = 32'h3000022c /* 0x02a0 */;
            169: data_o = 32'h30000224 /* 0x02a4 */;
            170: data_o = 32'h00000000 /* 0x02a8 */;
            171: data_o = 32'h00000000 /* 0x02ac */;
            172: data_o = 32'h00000000 /* 0x02b0 */;
            173: data_o = 32'h00000000 /* 0x02b4 */;
            174: data_o = 32'h00000000 /* 0x02b8 */;
            175: data_o = 32'h00000000 /* 0x02bc */;
            176: data_o = 32'h00000000 /* 0x02c0 */;
            177: data_o = 32'h00000000 /* 0x02c4 */;
            178: data_o = 32'h00000000 /* 0x02c8 */;
            179: data_o = 32'h00000000 /* 0x02cc */;
            180: data_o = 32'h00000000 /* 0x02d0 */;
            181: data_o = 32'h00000000 /* 0x02d4 */;
            182: data_o = 32'h00000000 /* 0x02d8 */;
            183: data_o = 32'h00000000 /* 0x02dc */;
            184: data_o = 32'h00000000 /* 0x02e0 */;
            185: data_o = 32'h00000000 /* 0x02e4 */;
            186: data_o = 32'h00000000 /* 0x02e8 */;
            187: data_o = 32'h00000000 /* 0x02ec */;
            188: data_o = 32'h00000000 /* 0x02f0 */;
            189: data_o = 32'h00000000 /* 0x02f4 */;
            190: data_o = 32'h00000000 /* 0x02f8 */;
            191: data_o = 32'h00000000 /* 0x02fc */;
            192: data_o = 32'h00000000 /* 0x0300 */;
            193: data_o = 32'h00000000 /* 0x0304 */;
            194: data_o = 32'h00000000 /* 0x0308 */;
            195: data_o = 32'h00000000 /* 0x030c */;
            196: data_o = 32'h00000000 /* 0x0310 */;
            197: data_o = 32'h00000000 /* 0x0314 */;
            198: data_o = 32'h00000000 /* 0x0318 */;
            199: data_o = 32'h00000000 /* 0x031c */;
            200: data_o = 32'h00000000 /* 0x0320 */;
            201: data_o = 32'h00000000 /* 0x0324 */;
            202: data_o = 32'h00000000 /* 0x0328 */;
            203: data_o = 32'h00000000 /* 0x032c */;
            204: data_o = 32'h00000000 /* 0x0330 */;
            205: data_o = 32'h00000000 /* 0x0334 */;
            206: data_o = 32'h00000000 /* 0x0338 */;
            207: data_o = 32'h00000000 /* 0x033c */;
            208: data_o = 32'h00000000 /* 0x0340 */;
            209: data_o = 32'h00000000 /* 0x0344 */;
            210: data_o = 32'h00000000 /* 0x0348 */;
            211: data_o = 32'h00000000 /* 0x034c */;
            212: data_o = 32'h00000000 /* 0x0350 */;
            213: data_o = 32'h00000000 /* 0x0354 */;
            214: data_o = 32'h00000000 /* 0x0358 */;
            215: data_o = 32'h00000000 /* 0x035c */;
            216: data_o = 32'h00000000 /* 0x0360 */;
            217: data_o = 32'h00000000 /* 0x0364 */;
            218: data_o = 32'h00000000 /* 0x0368 */;
            219: data_o = 32'h00000000 /* 0x036c */;
            220: data_o = 32'h00000000 /* 0x0370 */;
            221: data_o = 32'h00000000 /* 0x0374 */;
            222: data_o = 32'h00000000 /* 0x0378 */;
            223: data_o = 32'h00000000 /* 0x037c */;
            224: data_o = 32'h00000000 /* 0x0380 */;
            225: data_o = 32'h00000000 /* 0x0384 */;
            226: data_o = 32'h00000000 /* 0x0388 */;
            227: data_o = 32'h00000000 /* 0x038c */;
            228: data_o = 32'h00000000 /* 0x0390 */;
            229: data_o = 32'h00000000 /* 0x0394 */;
            230: data_o = 32'h00000000 /* 0x0398 */;
            231: data_o = 32'h00000000 /* 0x039c */;
            232: data_o = 32'h00000000 /* 0x03a0 */;
            233: data_o = 32'h00000000 /* 0x03a4 */;
            234: data_o = 32'h00000000 /* 0x03a8 */;
            235: data_o = 32'h00000000 /* 0x03ac */;
            236: data_o = 32'h00000000 /* 0x03b0 */;
            237: data_o = 32'h00000000 /* 0x03b4 */;
            238: data_o = 32'h00000000 /* 0x03b8 */;
            239: data_o = 32'h00000000 /* 0x03bc */;
            240: data_o = 32'h00000000 /* 0x03c0 */;
            241: data_o = 32'h00000000 /* 0x03c4 */;
            242: data_o = 32'h00000000 /* 0x03c8 */;
            243: data_o = 32'h00000000 /* 0x03cc */;
            244: data_o = 32'h00000000 /* 0x03d0 */;
            245: data_o = 32'h00000000 /* 0x03d4 */;
            246: data_o = 32'h00000000 /* 0x03d8 */;
            247: data_o = 32'h00000000 /* 0x03dc */;
            248: data_o = 32'h00000000 /* 0x03e0 */;
            249: data_o = 32'h00000000 /* 0x03e4 */;
            250: data_o = 32'h00000000 /* 0x03e8 */;
            251: data_o = 32'h00000000 /* 0x03ec */;
            252: data_o = 32'h00000000 /* 0x03f0 */;
            253: data_o = 32'h00000000 /* 0x03f4 */;
            254: data_o = 32'h00000000 /* 0x03f8 */;
            255: data_o = 32'h00000000 /* 0x03fc */;
            default: data_o = '0;
        endcase
    end

endmodule

// Copyright 2022 ETH Zurich and University of Bologna.
// Solderpad Hardware License, Version 0.51, see LICENSE for details.
// SPDX-License-Identifier: SHL-0.51
//
// Fabian Schuiki <fschuiki@iis.ee.ethz.ch>
// Florian Zaruba <zarubaf@iis.ee.ethz.ch>
// Stefan Mach <smach@iis.ee.ethz.ch>
// Thomas Benz <tbenz@iis.ee.ethz.ch>
// Paul Scheffler <paulsc@iis.ee.ethz.ch>
// Wolfgang Roenninger <wroennin@iis.ee.ethz.ch>
//
// AUTOMATICALLY GENERATED by gen_bootrom.py; edit the script instead.

module snitch_bootrom #(
    parameter int unsigned AddrWidth = 32,
    parameter int unsigned DataWidth = 32
)(
    input  logic                 clk_i,
    input  logic                 rst_ni,
    input  logic                 req_i,
    input  logic [AddrWidth-1:0] addr_i,
    output logic [DataWidth-1:0] data_o
);
    localparam unsigned NumWords = 64;
    logic [$clog2(NumWords)-1:0] word;

    assign word = addr_i / (DataWidth / 8);

    always_comb begin
        data_o = '0;
        unique case (word)
        000: data_o = 32'h30057073 /* 0x0000 */;
            001: data_o = 32'h00000293 /* 0x0004 */;
            002: data_o = 32'h00000313 /* 0x0008 */;
            003: data_o = 32'h00000393 /* 0x000c */;
            004: data_o = 32'h00000413 /* 0x0010 */;
            005: data_o = 32'h00000493 /* 0x0014 */;
            006: data_o = 32'h00000513 /* 0x0018 */;
            007: data_o = 32'h00000593 /* 0x001c */;
            008: data_o = 32'h00000613 /* 0x0020 */;
            009: data_o = 32'h00000693 /* 0x0024 */;
            010: data_o = 32'h00000713 /* 0x0028 */;
            011: data_o = 32'h00000793 /* 0x002c */;
            012: data_o = 32'h00000813 /* 0x0030 */;
            013: data_o = 32'h00000893 /* 0x0034 */;
            014: data_o = 32'h00000913 /* 0x0038 */;
            015: data_o = 32'h00000993 /* 0x003c */;
            016: data_o = 32'h00000a13 /* 0x0040 */;
            017: data_o = 32'h00000a93 /* 0x0044 */;
            018: data_o = 32'h00000b13 /* 0x0048 */;
            019: data_o = 32'h00000b93 /* 0x004c */;
            020: data_o = 32'h00000c13 /* 0x0050 */;
            021: data_o = 32'h00000c93 /* 0x0054 */;
            022: data_o = 32'h00000d13 /* 0x0058 */;
            023: data_o = 32'h00000d93 /* 0x005c */;
            024: data_o = 32'h00000e13 /* 0x0060 */;
            025: data_o = 32'h00000e93 /* 0x0064 */;
            026: data_o = 32'h00000f13 /* 0x0068 */;
            027: data_o = 32'h00000f93 /* 0x006c */;
            028: data_o = 32'h05c000ef /* 0x0070 */;
            029: data_o = 32'h00000297 /* 0x0074 */;
            030: data_o = 32'h03c28293 /* 0x0078 */;
            031: data_o = 32'h30529073 /* 0x007c */;
            032: data_o = 32'h10500073 /* 0x0080 */;
            033: data_o = 32'h00001297 /* 0x0084 */;
            034: data_o = 32'hf7c28293 /* 0x0088 */;
            035: data_o = 32'h0002a283 /* 0x008c */;
            036: data_o = 32'h000280e7 /* 0x0090 */;
            037: data_o = 32'h00001297 /* 0x0094 */;
            038: data_o = 32'hf6c28293 /* 0x0098 */;
            039: data_o = 32'h0052a223 /* 0x009c */;
            040: data_o = 32'hf61ff06f /* 0x00a0 */;
            041: data_o = 32'h00000013 /* 0x00a4 */;
            042: data_o = 32'h00000013 /* 0x00a8 */;
            043: data_o = 32'h00000013 /* 0x00ac */;
            044: data_o = 32'h02040fb7 /* 0x00b0 */;
            045: data_o = 32'h00000f13 /* 0x00b4 */;
            046: data_o = 32'h03efa423 /* 0x00b8 */;
            047: data_o = 32'h30200073 /* 0x00bc */;
            048: data_o = 32'h00008067 /* 0x00c0 */;
            049: data_o = 32'h00000000 /* 0x00c4 */;
            050: data_o = 32'h00000000 /* 0x00c8 */;
            051: data_o = 32'h304467f3 /* 0x00cc */;
            052: data_o = 32'h300467f3 /* 0x00d0 */;
            053: data_o = 32'h00008067 /* 0x00d4 */;
            054: data_o = 32'h00000000 /* 0x00d8 */;
            055: data_o = 32'h00000000 /* 0x00dc */;
            056: data_o = 32'h00000000 /* 0x00e0 */;
            057: data_o = 32'h00000000 /* 0x00e4 */;
            058: data_o = 32'h00000000 /* 0x00e8 */;
            059: data_o = 32'h00000000 /* 0x00ec */;
            060: data_o = 32'h00000000 /* 0x00f0 */;
            061: data_o = 32'h00000000 /* 0x00f4 */;
            062: data_o = 32'h00000000 /* 0x00f8 */;
            063: data_o = 32'h00000000 /* 0x00fc */;
            default: data_o = '0;
        endcase
    end

endmodule
